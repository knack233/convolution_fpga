module    mul_medium
(
    input signed[8:0]   mul_1 ,
    input signed[8:0]   mul_2 ,
    input signed[8:0]   mul_3 ,
    input signed[8:0]   mul_4 ,
    input signed[8:0]   mul_5 ,
    input signed[8:0]   mul_6 ,
    input signed[8:0]   mul_7 ,
    input signed[8:0]   mul_8 ,
    input signed[8:0]   mul_9 ,
    input signed[8:0]   mul_11,
    input signed[8:0]   mul_22,
    input signed[8:0]   mul_33,
    input signed[8:0]   mul_44,
    input signed[8:0]   mul_55,
    input signed[8:0]   mul_66,
    input signed[8:0]   mul_77,
    input signed[8:0]   mul_88,
    input signed[8:0]   mul_99,    
    output signed [15:0] mul_S
);












endmodule